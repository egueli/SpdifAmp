package constants is
  -- FPGA board frequency
  constant clock_frequency : real := 50.0e6;

end package;