library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity top is
  port (
    clk : in std_logic;
    rst : in std_logic;
    input : in std_logic;
    output : out std_logic
  );
end top; 

architecture str of top is

begin

end architecture;