library spdif_amp;
use spdif_amp.constants.all;

package sim_constants is
  constant clock_period : time := 1 sec / clock_frequency;
end package;